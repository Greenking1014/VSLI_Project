module RegisterFile ();
    
endmodule