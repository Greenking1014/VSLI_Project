module pcALU (

);
    
endmodule