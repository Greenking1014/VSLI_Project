module pcALU (
    ports
);
    
endmodule