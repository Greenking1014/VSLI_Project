module fpALU (
    ports
);
    
endmodule